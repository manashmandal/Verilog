
module test_mux;


endmodule
